LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY hazard_detection is
  -- IFID_REGISTER1 & 2 are placeholder names
  PORT( IDEX_REGISTER : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IFID_REGISTER1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        IFID_REGISTER2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
        STALL_REQUEST : OUT STD_LOGIC);
END hazard_detection;

ARCHITECTURE hazard_detection_arch of hazard_detection is
BEGIN
  STALL_REQUEST <= '1' WHEN (IDEX_REGISTER = IFID_REGISTER1 or IDEX_REGISTER = IFID_REGISTER2)
                       ELSE '0';
END hazard_detection_arch;
